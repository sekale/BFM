`ifndef DEFINESPKG_VH
`define DEFINESPKG_VH

package definesPkg;

parameter APB_ADDR_WIDTH = 32;
parameter APB_DATA_WIDTH = 32;

endpackage
`endif